module draw(x, y);
	input x,y;
	
	
	

endmodule